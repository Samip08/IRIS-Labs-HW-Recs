`timescale 1 ns / 1 ps

module uart_tb;
	reg clk;
	always #5 clk = (clk === 1'b0);  //100MHz

	reg [5:0] reset_cnt = 0;
	wire resetn = &reset_cnt;

	always @(posedge clk) begin
		reset_cnt <= reset_cnt + !resetn;
	end

	localparam ser_half_period = 53;
	event ser_sample;

	initial begin
		$dumpfile("uart_tb.vcd");
		$dumpvars(0, uart_tb);

		repeat (6) begin
			repeat (50000) @(posedge clk);
		end
		$finish;
	end


	wire ser_rx;
	wire ser_tx;

	wire flash_csb;
	wire flash_clk;
	wire flash_io0;
	wire flash_io1;
	wire flash_io2;
	wire flash_io3;

	rvsoc_wrapper #(
		.MEM_WORDS(256)
	) uut (
		.clk          (clk),
		.resetn       (resetn),
		.sensor_clk   (clk),    
		.ser_rx       (ser_rx),
		.ser_tx       (ser_tx),
		.flash_csb    (flash_csb),
		.flash_clk    (flash_clk),
		.flash_io0    (flash_io0),
		.flash_io1    (flash_io1),
		.flash_io2    (flash_io2),
		.flash_io3    (flash_io3)
	);
	spiflash spiflash (
		.csb(flash_csb),
		.clk(flash_clk),
		.io0(flash_io0),
		.io1(flash_io1),
		.io2(flash_io2),
		.io3(flash_io3)
	);

	reg [7:0] buffer;

	always begin
		@(negedge ser_tx);

		repeat (ser_half_period) @(posedge clk);
		-> ser_sample;

		repeat (8) begin
			repeat (ser_half_period) @(posedge clk);
			repeat (ser_half_period) @(posedge clk);
			buffer = {ser_tx, buffer[7:1]};
			-> ser_sample;
		end

		repeat (ser_half_period) @(posedge clk);
		repeat (ser_half_period) @(posedge clk);
		-> ser_sample;

		if (buffer < 32 || buffer >= 127)
			$display("Serial data: %d", buffer);
		else
			$display("Serial data: '%c'", buffer);
	end
endmodule
